library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package pkg_exp_tbl is
  component exp_tbl_31 is
    port (x : in  std_logic_vector(4 - 1 downto 0);
          y : out std_logic_vector(3 - 1 downto 0));
  end component;
  component exp_tbl_37 is
    port (x : in  std_logic_vector(6 - 1 downto 0);
          y : out std_logic_vector(14 - 1 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 23 bits) avec 36 bits en sortie
  component log_tbl_40 is
    port (x : in  std_logic_vector(3 downto 0);
          y : out std_logic_vector(35 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 20 bits) avec 39 bits en sortie
  component log_tbl_43 is
    port (x : in  std_logic_vector(3 downto 0);
          y : out std_logic_vector(38 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 17 bits) avec 42 bits en sortie
  component log_tbl_46 is
    port (x : in  std_logic_vector(3 downto 0);
          y : out std_logic_vector(41 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 14 bits) avec 45 bits en sortie
  component log_tbl_49 is
    port (x : in  std_logic_vector(3 downto 0);
          y : out std_logic_vector(44 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 11 bits) avec 48 bits en sortie
  component log_tbl_52 is
    port (x : in  std_logic_vector(3 downto 0);
          y : out std_logic_vector(47 downto 0));
  end component;
  -- tabule e ^ x - x - 1 avec 5 bits en entree, 1 en sortie
  -- le dernier bit de l'entree est le 8eme apres la virgule
  component exp_tbl_56 is
    port (x : in  std_logic_vector(4 downto 0);
          y : out std_logic_vector(0 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 8 bits) avec 51 bits en sortie
  component log_tbl_56 is
    port (x : in  std_logic_vector(4 downto 0);
          y : out std_logic_vector(50 downto 0));
  end component;
  -- tabule e ^ x - x - 1 avec 4 bits en entree, 3 en sortie
  -- le dernier bit de l'entree est le 5eme apres la virgule
  -- l'entree a en plus un bit de signe
  component exp_tbl_58 is
    port (x : in  std_logic_vector(4 downto 0);
          y : out std_logic_vector(2 downto 0));
  end component;
  -- tabule ln(e ^ x tronque a 5 bits) avec 55 bits en sortie
  component log_tbl_58 is
    port (x : in  std_logic_vector(4 downto 0);
          y : out std_logic_vector(54 downto 0));
  end component;
end package;

-- tables pour le composant exp_31
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity exp_tbl_31 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of exp_tbl_31 is
begin
  with x select
    y <= "000" when "0000",
         "000" when "0001",
         "000" when "0010",
         "000" when "0011",
         "000" when "0100",
         "000" when "0101",
         "001" when "0110",
         "001" when "0111",
         "001" when "1000",
         "001" when "1001",
         "010" when "1010",
         "010" when "1011",
         "010" when "1100",
         "011" when "1101",
         "011" when "1110",
         "100" when "1111",
         "---" when others;
end architecture;

-- tables pour le composant exp_37
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity exp_tbl_37 is
  port ( x : in  std_logic_vector(5 downto 0);
         y : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of exp_tbl_37 is
begin
  with x select
    y <= "00000000000000" when "000000",
         "00000000000100" when "000001",
         "00000000010000" when "000010",
         "00000000100100" when "000011",
         "00000001000000" when "000100",
         "00000001100100" when "000101",
         "00000010010000" when "000110",
         "00000011000100" when "000111",
         "00000100000000" when "001000",
         "00000101000100" when "001001",
         "00000110010000" when "001010",
         "00000111100100" when "001011",
         "00001001000000" when "001100",
         "00001010100100" when "001101",
         "00001100010000" when "001110",
         "00001110000100" when "001111",
         "00010000000000" when "010000",
         "00010010000100" when "010001",
         "00010100010000" when "010010",
         "00010110100100" when "010011",
         "00011001000000" when "010100",
         "00011011100100" when "010101",
         "00011110010000" when "010110",
         "00100001000100" when "010111",
         "00100100000000" when "011000",
         "00100111000100" when "011001",
         "00101010010000" when "011010",
         "00101101100100" when "011011",
         "00110001000000" when "011100",
         "00110100100100" when "011101",
         "00111000010000" when "011110",
         "00111100000100" when "011111",
         "01000000000000" when "100000",
         "01000100000100" when "100001",
         "01001000010000" when "100010",
         "01001100100100" when "100011",
         "01010001000000" when "100100",
         "01010101100100" when "100101",
         "01011010010000" when "100110",
         "01011111000100" when "100111",
         "01100100000000" when "101000",
         "01101001000100" when "101001",
         "01101110010000" when "101010",
         "01110011100100" when "101011",
         "01111001000000" when "101100",
         "01111110100100" when "101101",
         "10000100010000" when "101110",
         "10001010000100" when "101111",
         "10010000000000" when "110000",
         "10010110000100" when "110001",
         "10011100010000" when "110010",
         "10100010100100" when "110011",
         "10101001000000" when "110100",
         "10101111100100" when "110101",
         "10110110010000" when "110110",
         "10111101000100" when "110111",
         "11000100000000" when "111000",
         "11001011000100" when "111001",
         "11010010010000" when "111010",
         "11011001100100" when "111011",
         "11100001000000" when "111100",
         "11101000100100" when "111101",
         "11110000010000" when "111110",
         "11111000000100" when "111111",
         "--------------" when others;
end architecture;

-- tables pour le composant exp_40
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_40 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(35 downto 0) );
end entity;

architecture arch of log_tbl_40 is
begin
  with x select
    y <= "000000000000000000000000000000000000" when "0000",
         "000000000000000000000001000000000000" when "0001",
         "000000000000000000000100000000000000" when "0010",
         "000000000000000000001001000000000000" when "0011",
         "000000000000000000010000000000000000" when "0100",
         "000000000000000000011001000000000000" when "0101",
         "000000000000000000100100000000000000" when "0110",
         "000000000000000000110001000000000000" when "0111",
         "000000000000000001000000000000000000" when "1000",
         "000000000000000001010001000000000000" when "1001",
         "000000000000000001100100000000000000" when "1010",
         "000000000000000001111001000000000000" when "1011",
         "000000000000000010001111111111111111" when "1100",
         "000000000000000010101000111111111111" when "1101",
         "000000000000000011000011111111111111" when "1110",
         "000000000000000011100000111111111111" when "1111",
         "------------------------------------" when others;
end architecture;

-- tables pour le composant exp_43
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_43 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(38 downto 0) );
end entity;

architecture arch of log_tbl_43 is
begin
  with x select
    y <= "000000000000000000000000000000000000000" when "0000",
         "000000000000000000001000000000000000000" when "0001",
         "000000000000000000011111111111111111111" when "0010",
         "000000000000000001000111111111111111100" when "0011",
         "000000000000000001111111111111111110101" when "0100",
         "000000000000000011000111111111111101011" when "0101",
         "000000000000000100011111111111111011100" when "0110",
         "000000000000000110000111111111111000111" when "0111",
         "000000000000000111111111111111110101011" when "1000",
         "000000000000001010000111111111110000111" when "1001",
         "000000000000001100011111111111101011001" when "1010",
         "000000000000001111000111111111100100010" when "1011",
         "000000000000010001111111111111011100000" when "1100",
         "000000000000010101000111111111010010010" when "1101",
         "000000000000011000011111111111000110111" when "1110",
         "000000000000011100000111111110111001110" when "1111",
         "---------------------------------------" when others;
end architecture;

-- tables pour le composant exp_46
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_46 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(41 downto 0) );
end entity;

architecture arch of log_tbl_46 is
begin
  with x select
    y <= "000000000000000000000000000000000000000000" when "0000",
         "000000000000000000111111111111111110101011" when "0001",
         "000000000000000011111111111111110101010101" when "0010",
         "000000000000001000111111111111011100000000" when "0011",
         "000000000000001111111111111110101010101011" when "0100",
         "000000000000011000111111111101011001010110" when "0101",
         "000000000000100011111111111011100000000001" when "0110",
         "000000000000110000111111111000110110101100" when "0111",
         "000000000000111111111111110101010101010111" when "1000",
         "000000000001010000111111110000110100000011" when "1001",
         "000000000001100011111111101011001010110000" when "1010",
         "000000000001111000111111100100010001011100" when "1011",
         "000000000010001111111111011100000000001010" when "1100",
         "000000000010101000111111010010001110111001" when "1101",
         "000000000011000011111111000110110101101000" when "1110",
         "000000000011100000111110111001101100011001" when "1111",
         "------------------------------------------" when others;
end architecture;

-- tables pour le composant exp_49
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_49 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(44 downto 0) );
end entity;

architecture arch of log_tbl_49 is
begin
  with x select
    y <= "000000000000000000000000000000000000000000000" when "0000",
         "000000000000000111111111111110101010101010111" when "0001",
         "000000000000011111111111110101010101011001011" when "0010",
         "000000000001000111111111011100000000010100010" when "0011",
         "000000000001111111111110101010101011101010101" when "0100",
         "000000000011000111111101011001010111110001100" when "0101",
         "000000000100011111111011100000000101000011111" when "0110",
         "000000000110000111111000110110110100000010110" when "0111",
         "000000000111111111110101010101100101010100111" when "1000",
         "000000001010000111110000110100011001100111100" when "1001",
         "000000001100011111101011001011010001101101100" when "1010",
         "000000001111000111100100010010001110011111101" when "1011",
         "000000010001111111011100000001010000111101000" when "1100",
         "000000010101000111010010010000011010001010011" when "1101",
         "000000011000011111000110110111101011010010110" when "1110",
         "000000011100000110111001101111000101100111000" when "1111",
         "---------------------------------------------" when others;
end architecture;

-- tables pour le composant exp_52
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_52 is
  port ( x : in  std_logic_vector(3 downto 0);
         y : out std_logic_vector(47 downto 0) );
end entity;

architecture arch of log_tbl_52 is
begin
  with x select
    y <= "000000000000000000000000000000000000000000000000" when "0000",
         "000000000000111111111110101010101100101010100111" when "0001",
         "000000000011111111110101010101110101010011101111" when "0010",
         "000000001000111111011100000010100001110011110111" when "0011",
         "000000001111111110101010110010101001110111100011" when "0100",
         "000000011000111101011001101000110100111001011010" when "0101",
         "000000100011111011100000101000011001111100001001" when "0110",
         "000000110000111000110111110101011111100100101101" when "0111",
         "000000111111110101010111010100111011110100010000" when "1000",
         "000001010000110000110111001100010100000010010101" when "1001",
         "000001100011101011001111100001111100110110111011" when "1010",
         "000001111000100100011000011100111010000100101010" when "1011",
         "000010001111011100001010000100111110100010110110" when "1100",
         "000010101000010010011100100010101100000111101100" when "1101",
         "000011000011000111000111111111010011100010011100" when "1110",
         "000011011111111010000100100100110100010101100011" when "1111",
         "------------------------------------------------" when others;
end architecture;

-- tables pour le composant exp_56
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity exp_tbl_56 is
  port ( x : in  std_logic_vector(4 downto 0);
         y : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of exp_tbl_56 is
begin
  with x select
    y <= "0" when "00000",
         "0" when "00001",
         "0" when "00010",
         "0" when "00011",
         "0" when "00100",
         "0" when "00101",
         "0" when "00110",
         "0" when "00111",
         "0" when "01000",
         "0" when "01001",
         "0" when "01010",
         "0" when "01011",
         "0" when "01100",
         "0" when "01101",
         "0" when "01110",
         "0" when "01111",
         "0" when "10000",
         "0" when "10001",
         "0" when "10010",
         "0" when "10011",
         "0" when "10100",
         "0" when "10101",
         "0" when "10110",
         "1" when "10111",
         "1" when "11000",
         "1" when "11001",
         "1" when "11010",
         "1" when "11011",
         "1" when "11100",
         "1" when "11101",
         "1" when "11110",
         "1" when "11111",
         "-" when others;
end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_56 is
  port ( x : in  std_logic_vector(4 downto 0);
         y : out std_logic_vector(50 downto 0) );
end entity;

architecture arch of log_tbl_56 is
begin
  with x select
    y <= "000000000000000000000000000000000000000000000000000" when "00000",
         "000000000111111110101010111010100111011110100010000" when "00001",
         "000000011111110101011001010011101111100110000111100" when "00010",
         "000001000111011100010100000011111101111010110001001" when "00011",
         "000001111110101011101001111000000111111110000011100" when "00100",
         "000011000101011011101111001011100101011010100010110" when "00101",
         "000100011011100100111110000010101001001110111001011" when "00110",
         "000110000000111111110110000101000001101110011010000" when "00111",
         "000111110101100100111100011000011111001100111111111" when "01000",
         "001001111001001100111011011011100001001101000000001" when "01001",
         "001100001011110000100011000000001010000101010000001" when "01010",
         "001110101101001000101000000110111000110110010101110" when "01011",
         "010001011101001110000100111001101001000110000001111" when "01100",
         "010100011011111001111000100110111000111000001010010" when "01101",
         "010111101001000101000111011100110100011100100000101" when "01110",
         "011011000100101000111010100100100111101001010111000" when "01111",
         "011110101110011110011111111101110100111010101100110" when "10000",
         "100010100110011111001010011001110001101110001110110" when "10001",
         "100110101100100100010001010111001000010100011111001" when "10010",
         "101011000000100111010000111101011110101111101001000" when "10011",
         "101111100010100001101001111001000010111000101111011" when "10100",
         "110100010010001101000001010110011011100100001111110" when "10101",
         "111001001111100011000000111110011110011111000000101" when "10110",
         "000011110010110101110101000110101001010010110100011" when "10111",
         "001001011000100110010010100001001110110100110011100" when "11000",
         "001111001011101000101001110011100110010011011111000" when "11001",
         "010101001011110110111001110111111100110001010011001" when "11010",
         "011011011001001011000101101101010010101010011100101" when "11011",
         "100001110011011111010100010011110001001001011111000" when "11100",
         "101000011010101101110000101001000011100010111100111" when "11101",
         "101111001110110000101001100100110100110010100010101" when "11110",
         "110110001111100010010001110101010000110100011010001" when "11111",
         "---------------------------------------------------" when others;
end architecture;

-- tables pour le composant exp_58
-- ===============================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity exp_tbl_58 is
  port ( x : in  std_logic_vector(4 downto 0);
         y : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of exp_tbl_58 is
begin
  with x select
    y <= "011" when "11111",
         "011" when "11110",
         "010" when "11101",
         "010" when "11100",
         "001" when "11011",
         "001" when "11010",
         "001" when "11001",
         "001" when "11000",
         "000" when "10111",
         "000" when "10110",
         "000" when "10101",
         "000" when "10100",
         "000" when "10011",
         "000" when "10010",
         "000" when "10001",
         "000" when "10000",
         "000" when "00000",
         "000" when "00001",
         "000" when "00010",
         "000" when "00011",
         "000" when "00100",
         "000" when "00101",
         "000" when "00110",
         "000" when "00111",
         "001" when "01000",
         "001" when "01001",
         "001" when "01010",
         "010" when "01011",
         "010" when "01100",
         "011" when "01101",
         "011" when "01110",
         "100" when "01111",
         "---" when others;
end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity log_tbl_58 is
  port ( x : in  std_logic_vector(4 downto 0);
         y : out std_logic_vector(54 downto 0) );
end entity;

architecture arch of log_tbl_58 is
begin
  with x select
    y <= "0101011100111011011100010110100000101010011111010010001" when "11111",
         "0000010100100010100001101000100111001001101100110110011" when "11110",
         "1000010100100010100001101000100111001001101100110110011" when "11101",
         "0011110101001010010101001001001000110011011101000001101" when "11100",
         "1011110101001010010101001001001000110011011101000001101" when "11011",
         "0111111010111110100011101111011000000101010001101111110" when "11010",
         "0100100010101011100000011100111000101000111101011111010" when "11001",
         "0001101001011000100001000100110100110110111001001001111" when "11000",
         "1001101001011000100001000100110100110110111001001001111" when "10111",
         "0111001100100011100011011001011001110110011011110011000" when "10110",
         "0101001001111101101001111001000101011011001111000110111" when "10101",
         "0011011111101000000011010110101010000111101101100100000" when "10100",
         "0010001011110001110100000100010011111100100011110111110" when "10011",
         "0001001100110101111001011101010110010100100110001000101" when "10010",
         "0000100001011001100010110101100111100011101000000110100" when "10001",
         "0000001000001010111011000100111100111010001000100010010" when "10000",
         "0000000000000000000000000000000000000000000000000000000" when "00000",
         "0000000111110101100100111100011000011111001100111111111" when "00001",
         "0000011110101110011110011111111101110100111010101100110" when "00010",
         "0001000011110010110101110101000110101001010010110100011" when "00011",
         "0001110110001111100010010001110101010000110100011010001" when "00100",
         "0010110101010101101000001111110000000001010110111001011" when "00101",
         "0100000000011001111100011110101100001101100001011000011" when "00110",
         "0101010110110100101011000110000101110101001010010111001" when "00111",
         "0000100011011100111100100101010000111000001110101010111" when "01000",
         "0010011000101000110101010001010100010110011111001000000" when "01001",
         "0100010111000111010100010100011110111000101100111101100" when "01010",
         "0000101110010000100100000010100111111101100011010110110" when "01011",
         "0011000110001010000000100101000100001011111111100101100" when "01100",
         "0000001100110111000001001101000000011001111011010000010" when "01101",
         "0010111011000010001000010000110011011100001001110101110" when "01110",
         "0000101011100101011111101100111110001110110101111101000" when "01111",
         "-------------------------------------------------------" when others;
end architecture;

